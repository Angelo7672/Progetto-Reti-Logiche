-- test : sequenza di lunghezza massima, cio� RAM(0) = "11111111"

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity project_tb_seqmax is
end project_tb_seqmax;

architecture projecttb of project_tb_seqmax is
constant c_CLOCK_PERIOD         : time := 100 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);

signal RAM: ram_type := (
                        0 => std_logic_vector(to_unsigned( 255,8)),
			            1 => std_logic_vector(to_unsigned( 255,8)),
			            2 => std_logic_vector(to_unsigned( 222,8)),
			            3 => std_logic_vector(to_unsigned( 145,8)),
                        4 => std_logic_vector(to_unsigned( 250,8)),
                        5 => std_logic_vector(to_unsigned( 140,8)),
                        6 => std_logic_vector(to_unsigned( 74,8)),
                        7 => std_logic_vector(to_unsigned( 158,8)),
                        8 => std_logic_vector(to_unsigned( 180,8)),
                        9 => std_logic_vector(to_unsigned( 111,8)),
                        10 => std_logic_vector(to_unsigned( 182,8)),
                        11 => std_logic_vector(to_unsigned( 79,8)),
                        12 => std_logic_vector(to_unsigned( 239,8)),
                        13 => std_logic_vector(to_unsigned( 238,8)),
                        14 => std_logic_vector(to_unsigned( 219,8)),
                        15 => std_logic_vector(to_unsigned( 93,8)),
                        16 => std_logic_vector(to_unsigned( 26,8)),
                        17 => std_logic_vector(to_unsigned( 89,8)),
                        18 => std_logic_vector(to_unsigned( 11,8)),
                        19 => std_logic_vector(to_unsigned( 63,8)),
                        20 => std_logic_vector(to_unsigned( 255,8)),
                        21 => std_logic_vector(to_unsigned( 255,8)),
                        22 => std_logic_vector(to_unsigned( 253,8)),
                        23 => std_logic_vector(to_unsigned( 98,8)),
                        24 => std_logic_vector(to_unsigned( 228,8)),
                        25 => std_logic_vector(to_unsigned( 59,8)),
                        26 => std_logic_vector(to_unsigned( 170,8)),
                        27 => std_logic_vector(to_unsigned( 54,8)),
                        28 => std_logic_vector(to_unsigned( 27,8)),
                        29 => std_logic_vector(to_unsigned( 194,8)),
                        30 => std_logic_vector(to_unsigned( 117,8)),
                        31 => std_logic_vector(to_unsigned( 145,8)),
                        32 => std_logic_vector(to_unsigned( 102,8)),
                        33 => std_logic_vector(to_unsigned( 244,8)),
                        34 => std_logic_vector(to_unsigned( 240,8)),
                        35 => std_logic_vector(to_unsigned( 231,8)),
                        36 => std_logic_vector(to_unsigned( 220,8)),
                        37 => std_logic_vector(to_unsigned( 95,8)),
                        38 => std_logic_vector(to_unsigned( 243,8)),
                        39 => std_logic_vector(to_unsigned( 88,8)),
                        40 => std_logic_vector(to_unsigned( 128,8)),
                        41 => std_logic_vector(to_unsigned( 10,8)),
                        42 => std_logic_vector(to_unsigned( 161,8)),
                        43 => std_logic_vector(to_unsigned( 135,8)),
                        44 => std_logic_vector(to_unsigned( 175,8)),
                        45 => std_logic_vector(to_unsigned( 18,8)),
                        46 => std_logic_vector(to_unsigned( 140,8)),
                        47 => std_logic_vector(to_unsigned( 96,8)),
                        48 => std_logic_vector(to_unsigned( 53,8)),
                        49 => std_logic_vector(to_unsigned( 192,8)),
                        50 => std_logic_vector(to_unsigned( 123,8)),
                        51 => std_logic_vector(to_unsigned( 225,8)),
                        52 => std_logic_vector(to_unsigned( 197,8)),
                        53 => std_logic_vector(to_unsigned( 127,8)),
                        54 => std_logic_vector(to_unsigned( 42,8)),
                        55 => std_logic_vector(to_unsigned( 253,8)),
                        56 => std_logic_vector(to_unsigned( 88,8)),
                        57 => std_logic_vector(to_unsigned( 17,8)),
                        58 => std_logic_vector(to_unsigned( 118,8)),
                        59 => std_logic_vector(to_unsigned( 171,8)),
                        60 => std_logic_vector(to_unsigned( 232,8)),
                        61 => std_logic_vector(to_unsigned( 72,8)),
                        62 => std_logic_vector(to_unsigned( 51,8)),
                        63 => std_logic_vector(to_unsigned( 28,8)),
                        64 => std_logic_vector(to_unsigned( 221,8)),
                        65 => std_logic_vector(to_unsigned( 148,8)),
                        66 => std_logic_vector(to_unsigned( 205,8)),
                        67 => std_logic_vector(to_unsigned( 224,8)),
                        68 => std_logic_vector(to_unsigned( 188,8)),
                        69 => std_logic_vector(to_unsigned( 192,8)),
                        70 => std_logic_vector(to_unsigned( 36,8)),
                        71 => std_logic_vector(to_unsigned( 209,8)),
                        72 => std_logic_vector(to_unsigned( 55,8)),
                        73 => std_logic_vector(to_unsigned( 3,8)),
                        74 => std_logic_vector(to_unsigned( 101,8)),
                        75 => std_logic_vector(to_unsigned( 68,8)),
                        76 => std_logic_vector(to_unsigned( 113,8)),
                        77 => std_logic_vector(to_unsigned( 192,8)),
                        78 => std_logic_vector(to_unsigned( 164,8)),
                        79 => std_logic_vector(to_unsigned( 131,8)),
                        80 => std_logic_vector(to_unsigned( 35,8)),
                        81 => std_logic_vector(to_unsigned( 148,8)),
                        82 => std_logic_vector(to_unsigned( 16,8)),
                        83 => std_logic_vector(to_unsigned( 134,8)),
                        84 => std_logic_vector(to_unsigned( 135,8)),
                        85 => std_logic_vector(to_unsigned( 88,8)),
                        86 => std_logic_vector(to_unsigned( 138,8)),
                        87 => std_logic_vector(to_unsigned( 127,8)),
                        88 => std_logic_vector(to_unsigned( 140,8)),
                        89 => std_logic_vector(to_unsigned( 205,8)),
                        90 => std_logic_vector(to_unsigned( 37,8)),
                        91 => std_logic_vector(to_unsigned( 108,8)),
                        92 => std_logic_vector(to_unsigned( 67,8)),
                        93 => std_logic_vector(to_unsigned( 73,8)),
                        94 => std_logic_vector(to_unsigned( 59,8)),
                        95 => std_logic_vector(to_unsigned( 219,8)),
                        96 => std_logic_vector(to_unsigned( 198,8)),
                        97 => std_logic_vector(to_unsigned( 183,8)),
                        98 => std_logic_vector(to_unsigned( 107,8)),
                        99 => std_logic_vector(to_unsigned( 248,8)),
                        100 => std_logic_vector(to_unsigned( 158,8)),
                        101 => std_logic_vector(to_unsigned( 130,8)),
                        102 => std_logic_vector(to_unsigned( 184,8)),
                        103 => std_logic_vector(to_unsigned( 50,8)),
                        104 => std_logic_vector(to_unsigned( 54,8)),
                        105 => std_logic_vector(to_unsigned( 181,8)),
                        106 => std_logic_vector(to_unsigned( 7,8)),
                        107 => std_logic_vector(to_unsigned( 44,8)),
                        108 => std_logic_vector(to_unsigned( 66,8)),
                        109 => std_logic_vector(to_unsigned( 61,8)),
                        110 => std_logic_vector(to_unsigned( 200,8)),
                        111 => std_logic_vector(to_unsigned( 150,8)),
                        112 => std_logic_vector(to_unsigned( 163,8)),
                        113 => std_logic_vector(to_unsigned( 180,8)),
                        114 => std_logic_vector(to_unsigned( 32,8)),
                        115 => std_logic_vector(to_unsigned( 226,8)),
                        116 => std_logic_vector(to_unsigned( 89,8)),
                        117 => std_logic_vector(to_unsigned( 120,8)),
                        118 => std_logic_vector(to_unsigned( 80,8)),
                        119 => std_logic_vector(to_unsigned( 189,8)),
                        120 => std_logic_vector(to_unsigned( 27,8)),
                        121 => std_logic_vector(to_unsigned( 59,8)),
                        122 => std_logic_vector(to_unsigned( 186,8)),
                        123 => std_logic_vector(to_unsigned( 206,8)),
                        124 => std_logic_vector(to_unsigned( 194,8)),
                        125 => std_logic_vector(to_unsigned( 153,8)),
                        126 => std_logic_vector(to_unsigned( 95,8)),
                        127 => std_logic_vector(to_unsigned( 189,8)),
                        128 => std_logic_vector(to_unsigned( 215,8)),
                        129 => std_logic_vector(to_unsigned( 12,8)),
                        130 => std_logic_vector(to_unsigned( 22,8)),
                        131 => std_logic_vector(to_unsigned( 241,8)),
                        132 => std_logic_vector(to_unsigned( 66,8)),
                        133 => std_logic_vector(to_unsigned( 149,8)),
                        134 => std_logic_vector(to_unsigned( 204,8)),
                        135 => std_logic_vector(to_unsigned( 230,8)),
                        136 => std_logic_vector(to_unsigned( 172,8)),
                        137 => std_logic_vector(to_unsigned( 84,8)),
                        138 => std_logic_vector(to_unsigned( 222,8)),
                        139 => std_logic_vector(to_unsigned( 216,8)),
                        140 => std_logic_vector(to_unsigned( 141,8)),
                        141 => std_logic_vector(to_unsigned( 17,8)),
                        142 => std_logic_vector(to_unsigned( 239,8)),
                        143 => std_logic_vector(to_unsigned( 49,8)),
                        144 => std_logic_vector(to_unsigned( 214,8)),
                        145 => std_logic_vector(to_unsigned( 40,8)),
                        146 => std_logic_vector(to_unsigned( 98,8)),
                        147 => std_logic_vector(to_unsigned( 172,8)),
                        148 => std_logic_vector(to_unsigned( 145,8)),
                        149 => std_logic_vector(to_unsigned( 156,8)),
                        150 => std_logic_vector(to_unsigned( 47,8)),
                        151 => std_logic_vector(to_unsigned( 98,8)),
                        152 => std_logic_vector(to_unsigned( 37,8)),
                        153 => std_logic_vector(to_unsigned( 124,8)),
                        154 => std_logic_vector(to_unsigned( 48,8)),
                        155 => std_logic_vector(to_unsigned( 251,8)),
                        156 => std_logic_vector(to_unsigned( 235,8)),
                        157 => std_logic_vector(to_unsigned( 12,8)),
                        158 => std_logic_vector(to_unsigned( 49,8)),
                        159 => std_logic_vector(to_unsigned( 210,8)),
                        160 => std_logic_vector(to_unsigned( 92,8)),
                        161 => std_logic_vector(to_unsigned( 39,8)),
                        162 => std_logic_vector(to_unsigned( 63,8)),
                        163 => std_logic_vector(to_unsigned( 109,8)),
                        164 => std_logic_vector(to_unsigned( 237,8)),
                        165 => std_logic_vector(to_unsigned( 155,8)),
                        166 => std_logic_vector(to_unsigned( 136,8)),
                        167 => std_logic_vector(to_unsigned( 178,8)),
                        168 => std_logic_vector(to_unsigned( 132,8)),
                        169 => std_logic_vector(to_unsigned( 49,8)),
                        170 => std_logic_vector(to_unsigned( 71,8)),
                        171 => std_logic_vector(to_unsigned( 216,8)),
                        172 => std_logic_vector(to_unsigned( 199,8)),
                        173 => std_logic_vector(to_unsigned( 187,8)),
                        174 => std_logic_vector(to_unsigned( 59,8)),
                        175 => std_logic_vector(to_unsigned( 74,8)),
                        176 => std_logic_vector(to_unsigned( 1,8)),
                        177 => std_logic_vector(to_unsigned( 179,8)),
                        178 => std_logic_vector(to_unsigned( 164,8)),
                        179 => std_logic_vector(to_unsigned( 231,8)),
                        180 => std_logic_vector(to_unsigned( 93,8)),
                        181 => std_logic_vector(to_unsigned( 245,8)),
                        182 => std_logic_vector(to_unsigned( 31,8)),
                        183 => std_logic_vector(to_unsigned( 193,8)),
                        184 => std_logic_vector(to_unsigned( 113,8)),
                        185 => std_logic_vector(to_unsigned( 242,8)),
                        186 => std_logic_vector(to_unsigned( 0,8)),
                        187 => std_logic_vector(to_unsigned( 36,8)),
                        188 => std_logic_vector(to_unsigned( 231,8)),
                        189 => std_logic_vector(to_unsigned( 209,8)),
                        190 => std_logic_vector(to_unsigned( 218,8)),
                        191 => std_logic_vector(to_unsigned( 48,8)),
                        192 => std_logic_vector(to_unsigned( 125,8)),
                        193 => std_logic_vector(to_unsigned( 21,8)),
                        194 => std_logic_vector(to_unsigned( 92,8)),
                        195 => std_logic_vector(to_unsigned( 205,8)),
                        196 => std_logic_vector(to_unsigned( 122,8)),
                        197 => std_logic_vector(to_unsigned( 20,8)),
                        198 => std_logic_vector(to_unsigned( 129,8)),
                        199 => std_logic_vector(to_unsigned( 82,8)),
                        200 => std_logic_vector(to_unsigned( 76,8)),
                        201 => std_logic_vector(to_unsigned( 168,8)),
                        202 => std_logic_vector(to_unsigned( 235,8)),
                        203 => std_logic_vector(to_unsigned( 238,8)),
                        204 => std_logic_vector(to_unsigned( 215,8)),
                        205 => std_logic_vector(to_unsigned( 53,8)),
                        206 => std_logic_vector(to_unsigned( 212,8)),
                        207 => std_logic_vector(to_unsigned( 120,8)),
                        208 => std_logic_vector(to_unsigned( 251,8)),
                        209 => std_logic_vector(to_unsigned( 114,8)),
                        210 => std_logic_vector(to_unsigned( 250,8)),
                        211 => std_logic_vector(to_unsigned( 13,8)),
                        212 => std_logic_vector(to_unsigned( 125,8)),
                        213 => std_logic_vector(to_unsigned( 201,8)),
                        214 => std_logic_vector(to_unsigned( 56,8)),
                        215 => std_logic_vector(to_unsigned( 235,8)),
                        216 => std_logic_vector(to_unsigned( 149,8)),
                        217 => std_logic_vector(to_unsigned( 96,8)),
                        218 => std_logic_vector(to_unsigned( 142,8)),
                        219 => std_logic_vector(to_unsigned( 76,8)),
                        220 => std_logic_vector(to_unsigned( 114,8)),
                        221 => std_logic_vector(to_unsigned( 182,8)),
                        222 => std_logic_vector(to_unsigned( 209,8)),
                        223 => std_logic_vector(to_unsigned( 128,8)),
                        224 => std_logic_vector(to_unsigned( 117,8)),
                        225 => std_logic_vector(to_unsigned( 154,8)),
                        226 => std_logic_vector(to_unsigned( 28,8)),
                        227 => std_logic_vector(to_unsigned( 225,8)),
                        228 => std_logic_vector(to_unsigned( 35,8)),
                        229 => std_logic_vector(to_unsigned( 10,8)),
                        230 => std_logic_vector(to_unsigned( 59,8)),
                        231 => std_logic_vector(to_unsigned( 107,8)),
                        232 => std_logic_vector(to_unsigned( 245,8)),
                        233 => std_logic_vector(to_unsigned( 22,8)),
                        234 => std_logic_vector(to_unsigned( 126,8)),
                        235 => std_logic_vector(to_unsigned( 185,8)),
                        236 => std_logic_vector(to_unsigned( 12,8)),
                        237 => std_logic_vector(to_unsigned( 170,8)),
                        238 => std_logic_vector(to_unsigned( 131,8)),
                        239 => std_logic_vector(to_unsigned( 93,8)),
                        240 => std_logic_vector(to_unsigned( 112,8)),
                        241 => std_logic_vector(to_unsigned( 137,8)),
                        242 => std_logic_vector(to_unsigned( 186,8)),
                        243 => std_logic_vector(to_unsigned( 70,8)),
                        244 => std_logic_vector(to_unsigned( 247,8)),
                        245 => std_logic_vector(to_unsigned( 35,8)),
                        246 => std_logic_vector(to_unsigned( 31,8)),
                        247 => std_logic_vector(to_unsigned( 119,8)),
                        248 => std_logic_vector(to_unsigned( 160,8)),
                        249 => std_logic_vector(to_unsigned( 35,8)),
                        250 => std_logic_vector(to_unsigned( 64,8)),
                        251 => std_logic_vector(to_unsigned( 170,8)),
                        252 => std_logic_vector(to_unsigned( 197,8)),
                        253 => std_logic_vector(to_unsigned( 53,8)),
                        254 => std_logic_vector(to_unsigned( 178,8)),
                        255 => std_logic_vector(to_unsigned( 216,8)),
                        others => (others =>'0')); 
                         
component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;
                         
begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;

MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 2 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 2 ns;
            end if;
        end if;
    end if;
end process;

test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
    
    assert RAM(1000) = STD_LOGIC_VECTOR(TO_UNSIGNED(229, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1001) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1002) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1003) = STD_LOGIC_VECTOR(TO_UNSIGNED(150, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1004) = STD_LOGIC_VECTOR(TO_UNSIGNED(31, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1005) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1006) = STD_LOGIC_VECTOR(TO_UNSIGNED(149, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1007) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1008) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1009) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1010) = STD_LOGIC_VECTOR(TO_UNSIGNED(55, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1011) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1012) = STD_LOGIC_VECTOR(TO_UNSIGNED(31, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1013) = STD_LOGIC_VECTOR(TO_UNSIGNED(150, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1014) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1015) = STD_LOGIC_VECTOR(TO_UNSIGNED(135, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1016) = STD_LOGIC_VECTOR(TO_UNSIGNED(58, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1017) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1018) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1019) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1020) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1021) = STD_LOGIC_VECTOR(TO_UNSIGNED(229, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1022) = STD_LOGIC_VECTOR(TO_UNSIGNED(86, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1023) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1024) = STD_LOGIC_VECTOR(TO_UNSIGNED(86, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1025) = STD_LOGIC_VECTOR(TO_UNSIGNED(38, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1026) = STD_LOGIC_VECTOR(TO_UNSIGNED(40, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1027) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1028) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1029) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1030) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1031) = STD_LOGIC_VECTOR(TO_UNSIGNED(161, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1032) = STD_LOGIC_VECTOR(TO_UNSIGNED(244, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1033) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1034) = STD_LOGIC_VECTOR(TO_UNSIGNED(112, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1035) = STD_LOGIC_VECTOR(TO_UNSIGNED(210, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1036) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1037) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1038) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1039) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1040) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1041) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1042) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1043) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1044) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1045) = STD_LOGIC_VECTOR(TO_UNSIGNED(205, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1046) = STD_LOGIC_VECTOR(TO_UNSIGNED(38, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1047) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1048) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1049) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1050) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1051) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1052) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1053) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1054) = STD_LOGIC_VECTOR(TO_UNSIGNED(195, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1055) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1056) = STD_LOGIC_VECTOR(TO_UNSIGNED(91, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1057) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1058) = STD_LOGIC_VECTOR(TO_UNSIGNED(249, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1059) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1060) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1061) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1062) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1063) = STD_LOGIC_VECTOR(TO_UNSIGNED(250, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1064) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1065) = STD_LOGIC_VECTOR(TO_UNSIGNED(135, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1066) = STD_LOGIC_VECTOR(TO_UNSIGNED(229, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1067) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1068) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1069) = STD_LOGIC_VECTOR(TO_UNSIGNED(249, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1070) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1071) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1072) = STD_LOGIC_VECTOR(TO_UNSIGNED(52, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1073) = STD_LOGIC_VECTOR(TO_UNSIGNED(149, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1074) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1075) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1076) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1077) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1078) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1079) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1080) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1081) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1082) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1083) = STD_LOGIC_VECTOR(TO_UNSIGNED(195, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1084) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1085) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1086) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1087) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1088) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1089) = STD_LOGIC_VECTOR(TO_UNSIGNED(125, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1090) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1091) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1092) = STD_LOGIC_VECTOR(TO_UNSIGNED(58, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1093) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1094) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1095) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1096) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1097) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1098) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1099) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    
    assert RAM(1100) = STD_LOGIC_VECTOR(TO_UNSIGNED(86, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1101) = STD_LOGIC_VECTOR(TO_UNSIGNED(195, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1102) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1103) = STD_LOGIC_VECTOR(TO_UNSIGNED(52, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1104) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1105) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1106) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1107) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1108) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1109) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1110) = STD_LOGIC_VECTOR(TO_UNSIGNED(68, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1111) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1112) = STD_LOGIC_VECTOR(TO_UNSIGNED(3, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1113) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1114) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1115) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1116) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1117) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1118) = STD_LOGIC_VECTOR(TO_UNSIGNED(86, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1119) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1120) = STD_LOGIC_VECTOR(TO_UNSIGNED(55, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1121) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1122) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1123) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1124) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1125) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1126) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1127) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1128) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1129) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1130) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1131) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1132) = STD_LOGIC_VECTOR(TO_UNSIGNED(150, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1133) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1134) = STD_LOGIC_VECTOR(TO_UNSIGNED(210, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1135) = STD_LOGIC_VECTOR(TO_UNSIGNED(91, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1136) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1137) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1138) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1139) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1140) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1141) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1142) = STD_LOGIC_VECTOR(TO_UNSIGNED(126, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1143) = STD_LOGIC_VECTOR(TO_UNSIGNED(137, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1144) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1145) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1146) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1147) = STD_LOGIC_VECTOR(TO_UNSIGNED(244, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1148) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1149) = STD_LOGIC_VECTOR(TO_UNSIGNED(55, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1150) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1151) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1152) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1153) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1154) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1155) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1156) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1157) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1158) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1159) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1160) = STD_LOGIC_VECTOR(TO_UNSIGNED(111, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1161) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1162) = STD_LOGIC_VECTOR(TO_UNSIGNED(3, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1163) = STD_LOGIC_VECTOR(TO_UNSIGNED(112, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1164) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1165) = STD_LOGIC_VECTOR(TO_UNSIGNED(58, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1166) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1167) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1168) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1169) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1170) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1171) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1172) = STD_LOGIC_VECTOR(TO_UNSIGNED(249, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1173) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1174) = STD_LOGIC_VECTOR(TO_UNSIGNED(108, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1175) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1176) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1177) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1178) = STD_LOGIC_VECTOR(TO_UNSIGNED(125, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1179) = STD_LOGIC_VECTOR(TO_UNSIGNED(244, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1180) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1181) = STD_LOGIC_VECTOR(TO_UNSIGNED(43, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1182) = STD_LOGIC_VECTOR(TO_UNSIGNED(55, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1183) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1184) = STD_LOGIC_VECTOR(TO_UNSIGNED(135, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1185) = STD_LOGIC_VECTOR(TO_UNSIGNED(223, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1186) = STD_LOGIC_VECTOR(TO_UNSIGNED(126, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1187) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1188) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1189) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1190) = STD_LOGIC_VECTOR(TO_UNSIGNED(91, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1191) = STD_LOGIC_VECTOR(TO_UNSIGNED(58, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1192) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1193) = STD_LOGIC_VECTOR(TO_UNSIGNED(137, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1194) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1195) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1196) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1197) = STD_LOGIC_VECTOR(TO_UNSIGNED(108, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1198) = STD_LOGIC_VECTOR(TO_UNSIGNED(223, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1199) = STD_LOGIC_VECTOR(TO_UNSIGNED(150, 8)) report "TEST FALLITO" severity failure;
    
    assert RAM(1200) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1201) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1202) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1203) = STD_LOGIC_VECTOR(TO_UNSIGNED(108, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1204) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1205) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1206) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1207) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1208) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1209) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1210) = STD_LOGIC_VECTOR(TO_UNSIGNED(112, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1211) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1212) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1213) = STD_LOGIC_VECTOR(TO_UNSIGNED(43, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1214) = STD_LOGIC_VECTOR(TO_UNSIGNED(55, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1215) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1216) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1217) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1218) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1219) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1220) = STD_LOGIC_VECTOR(TO_UNSIGNED(223, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1221) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1222) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1223) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1224) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1225) = STD_LOGIC_VECTOR(TO_UNSIGNED(135, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1226) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1227) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1228) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1229) = STD_LOGIC_VECTOR(TO_UNSIGNED(205, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1230) = STD_LOGIC_VECTOR(TO_UNSIGNED(244, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1231) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1232) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1233) = STD_LOGIC_VECTOR(TO_UNSIGNED(108, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1234) = STD_LOGIC_VECTOR(TO_UNSIGNED(52, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1235) = STD_LOGIC_VECTOR(TO_UNSIGNED(112, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1236) = STD_LOGIC_VECTOR(TO_UNSIGNED(210, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1237) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1238) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1239) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1240) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1241) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1242) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1243) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1244) = STD_LOGIC_VECTOR(TO_UNSIGNED(43, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1245) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1246) = STD_LOGIC_VECTOR(TO_UNSIGNED(43, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1247) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1248) = STD_LOGIC_VECTOR(TO_UNSIGNED(31, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1249) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1250) = STD_LOGIC_VECTOR(TO_UNSIGNED(68, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1251) = STD_LOGIC_VECTOR(TO_UNSIGNED(149, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1252) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1253) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1254) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1255) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1256) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1257) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1258) = STD_LOGIC_VECTOR(TO_UNSIGNED(3, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1259) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1260) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1261) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1262) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1263) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1264) = STD_LOGIC_VECTOR(TO_UNSIGNED(31, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1265) = STD_LOGIC_VECTOR(TO_UNSIGNED(68, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1266) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1267) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1268) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1269) = STD_LOGIC_VECTOR(TO_UNSIGNED(250, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1270) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1271) = STD_LOGIC_VECTOR(TO_UNSIGNED(43, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1272) = STD_LOGIC_VECTOR(TO_UNSIGNED(52, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1273) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1274) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1275) = STD_LOGIC_VECTOR(TO_UNSIGNED(150, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1276) = STD_LOGIC_VECTOR(TO_UNSIGNED(40, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1277) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1278) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1279) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1280) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1281) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1282) = STD_LOGIC_VECTOR(TO_UNSIGNED(150, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1283) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1284) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1285) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1286) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1287) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1288) = STD_LOGIC_VECTOR(TO_UNSIGNED(205, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1289) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1290) = STD_LOGIC_VECTOR(TO_UNSIGNED(58, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1291) = STD_LOGIC_VECTOR(TO_UNSIGNED(205, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1292) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1293) = STD_LOGIC_VECTOR(TO_UNSIGNED(43, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1294) = STD_LOGIC_VECTOR(TO_UNSIGNED(223, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1295) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1296) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1297) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1298) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1299) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    
    assert RAM(1300) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1301) = STD_LOGIC_VECTOR(TO_UNSIGNED(205, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1302) = STD_LOGIC_VECTOR(TO_UNSIGNED(205, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1303) = STD_LOGIC_VECTOR(TO_UNSIGNED(244, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1304) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1305) = STD_LOGIC_VECTOR(TO_UNSIGNED(91, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1306) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1307) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1308) = STD_LOGIC_VECTOR(TO_UNSIGNED(229, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1309) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1310) = STD_LOGIC_VECTOR(TO_UNSIGNED(86, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1311) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1312) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1313) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1314) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1315) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1316) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1317) = STD_LOGIC_VECTOR(TO_UNSIGNED(125, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1318) = STD_LOGIC_VECTOR(TO_UNSIGNED(244, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1319) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1320) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1321) = STD_LOGIC_VECTOR(TO_UNSIGNED(249, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1322) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1323) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1324) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1325) = STD_LOGIC_VECTOR(TO_UNSIGNED(40, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1326) = STD_LOGIC_VECTOR(TO_UNSIGNED(150, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1327) = STD_LOGIC_VECTOR(TO_UNSIGNED(40, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1328) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1329) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1330) = STD_LOGIC_VECTOR(TO_UNSIGNED(108, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1331) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1332) = STD_LOGIC_VECTOR(TO_UNSIGNED(210, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1333) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1334) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1335) = STD_LOGIC_VECTOR(TO_UNSIGNED(55, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1336) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1337) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1338) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1339) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1340) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1341) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1342) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1343) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1344) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1345) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1346) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1347) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1348) = STD_LOGIC_VECTOR(TO_UNSIGNED(135, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1349) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1350) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1351) = STD_LOGIC_VECTOR(TO_UNSIGNED(3, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1352) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1353) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1354) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1355) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1356) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1357) = STD_LOGIC_VECTOR(TO_UNSIGNED(249, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1358) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1359) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1360) = STD_LOGIC_VECTOR(TO_UNSIGNED(149, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1361) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1362) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1363) = STD_LOGIC_VECTOR(TO_UNSIGNED(149, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1364) = STD_LOGIC_VECTOR(TO_UNSIGNED(91, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1365) = STD_LOGIC_VECTOR(TO_UNSIGNED(3, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1366) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1367) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1368) = STD_LOGIC_VECTOR(TO_UNSIGNED(149, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1369) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1370) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1371) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1372) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1373) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1374) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1375) = STD_LOGIC_VECTOR(TO_UNSIGNED(249, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1376) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1377) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1378) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1379) = STD_LOGIC_VECTOR(TO_UNSIGNED(161, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1380) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1381) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1382) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1383) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1384) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1385) = STD_LOGIC_VECTOR(TO_UNSIGNED(68, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1386) = STD_LOGIC_VECTOR(TO_UNSIGNED(68, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1387) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1388) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1389) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1390) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1391) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1392) = STD_LOGIC_VECTOR(TO_UNSIGNED(195, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1393) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1394) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1395) = STD_LOGIC_VECTOR(TO_UNSIGNED(3, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1396) = STD_LOGIC_VECTOR(TO_UNSIGNED(68, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1397) = STD_LOGIC_VECTOR(TO_UNSIGNED(125, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1398) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1399) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
   
    assert RAM(1400) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1401) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1402) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1403) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1404) = STD_LOGIC_VECTOR(TO_UNSIGNED(86, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1405) = STD_LOGIC_VECTOR(TO_UNSIGNED(38, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1406) = STD_LOGIC_VECTOR(TO_UNSIGNED(40, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1407) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1408) = STD_LOGIC_VECTOR(TO_UNSIGNED(190, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1409) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1410) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1411) = STD_LOGIC_VECTOR(TO_UNSIGNED(71, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1412) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1413) = STD_LOGIC_VECTOR(TO_UNSIGNED(108, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1414) = STD_LOGIC_VECTOR(TO_UNSIGNED(229, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1415) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1416) = STD_LOGIC_VECTOR(TO_UNSIGNED(137, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1417) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1418) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1419) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1420) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1421) = STD_LOGIC_VECTOR(TO_UNSIGNED(232, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1422) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1423) = STD_LOGIC_VECTOR(TO_UNSIGNED(88, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1424) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1425) = STD_LOGIC_VECTOR(TO_UNSIGNED(223, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1426) = STD_LOGIC_VECTOR(TO_UNSIGNED(126, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1427) = STD_LOGIC_VECTOR(TO_UNSIGNED(108, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1428) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1429) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1430) = STD_LOGIC_VECTOR(TO_UNSIGNED(111, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1431) = STD_LOGIC_VECTOR(TO_UNSIGNED(68, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1432) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1433) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1434) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1435) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1436) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1437) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1438) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1439) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1440) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1441) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1442) = STD_LOGIC_VECTOR(TO_UNSIGNED(40, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1443) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1444) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1445) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1446) = STD_LOGIC_VECTOR(TO_UNSIGNED(57, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1447) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1448) = STD_LOGIC_VECTOR(TO_UNSIGNED(175, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1449) = STD_LOGIC_VECTOR(TO_UNSIGNED(161, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1450) = STD_LOGIC_VECTOR(TO_UNSIGNED(195, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1451) = STD_LOGIC_VECTOR(TO_UNSIGNED(155, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1452) = STD_LOGIC_VECTOR(TO_UNSIGNED(230, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1453) = STD_LOGIC_VECTOR(TO_UNSIGNED(195, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1454) = STD_LOGIC_VECTOR(TO_UNSIGNED(125, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1455) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1456) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1457) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1458) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1459) = STD_LOGIC_VECTOR(TO_UNSIGNED(98, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1460) = STD_LOGIC_VECTOR(TO_UNSIGNED(138, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1461) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1462) = STD_LOGIC_VECTOR(TO_UNSIGNED(85, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1463) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1464) = STD_LOGIC_VECTOR(TO_UNSIGNED(115, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1465) = STD_LOGIC_VECTOR(TO_UNSIGNED(74, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1466) = STD_LOGIC_VECTOR(TO_UNSIGNED(249, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1467) = STD_LOGIC_VECTOR(TO_UNSIGNED(86, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1468) = STD_LOGIC_VECTOR(TO_UNSIGNED(18, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1469) = STD_LOGIC_VECTOR(TO_UNSIGNED(111, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1470) = STD_LOGIC_VECTOR(TO_UNSIGNED(112, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1471) = STD_LOGIC_VECTOR(TO_UNSIGNED(235, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1472) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1473) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1474) = STD_LOGIC_VECTOR(TO_UNSIGNED(28, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1475) = STD_LOGIC_VECTOR(TO_UNSIGNED(14, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1476) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1477) = STD_LOGIC_VECTOR(TO_UNSIGNED(152, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1478) = STD_LOGIC_VECTOR(TO_UNSIGNED(73, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1479) = STD_LOGIC_VECTOR(TO_UNSIGNED(176, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1480) = STD_LOGIC_VECTOR(TO_UNSIGNED(220, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1481) = STD_LOGIC_VECTOR(TO_UNSIGNED(223, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1482) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1483) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1484) = STD_LOGIC_VECTOR(TO_UNSIGNED(247, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1485) = STD_LOGIC_VECTOR(TO_UNSIGNED(58, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1486) = STD_LOGIC_VECTOR(TO_UNSIGNED(37, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1487) = STD_LOGIC_VECTOR(TO_UNSIGNED(137, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1488) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1489) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1490) = STD_LOGIC_VECTOR(TO_UNSIGNED(179, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1491) = STD_LOGIC_VECTOR(TO_UNSIGNED(149, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1492) = STD_LOGIC_VECTOR(TO_UNSIGNED(137, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1493) = STD_LOGIC_VECTOR(TO_UNSIGNED(137, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1494) = STD_LOGIC_VECTOR(TO_UNSIGNED(97, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1495) = STD_LOGIC_VECTOR(TO_UNSIGNED(192, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1496) = STD_LOGIC_VECTOR(TO_UNSIGNED(13, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1497) = STD_LOGIC_VECTOR(TO_UNSIGNED(206, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1498) = STD_LOGIC_VECTOR(TO_UNSIGNED(135, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1499) = STD_LOGIC_VECTOR(TO_UNSIGNED(0, 8)) report "TEST FALLITO" severity failure;
    
    assert RAM(1500) = STD_LOGIC_VECTOR(TO_UNSIGNED(209, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1501) = STD_LOGIC_VECTOR(TO_UNSIGNED(17, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1502) = STD_LOGIC_VECTOR(TO_UNSIGNED(43, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1503) = STD_LOGIC_VECTOR(TO_UNSIGNED(52, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1504) = STD_LOGIC_VECTOR(TO_UNSIGNED(126, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1505) = STD_LOGIC_VECTOR(TO_UNSIGNED(132, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1506) = STD_LOGIC_VECTOR(TO_UNSIGNED(162, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1507) = STD_LOGIC_VECTOR(TO_UNSIGNED(189, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1508) = STD_LOGIC_VECTOR(TO_UNSIGNED(40, 8)) report "TEST FALLITO" severity failure;
    assert RAM(1509) = STD_LOGIC_VECTOR(TO_UNSIGNED(172, 8)) report "TEST FALLITO" severity failure;
    
    assert false report "Simulation Ended! TEST PASSATO" severity failure;

end process test;    

end projecttb;

